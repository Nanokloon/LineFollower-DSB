module motorcontrol 
   (input logic clk,
    input logic reset,
    input logic direction, 
    input logic [?:0] count_in,
    output logic pwm);



endmodule
