module inputbuffer
   (input logic clk,
    input logic sensor_l_in,
    input logic sensor_m_in, 
    input logic sensor_r_in,
    output logic sensor_l_out,
    output logic sensor_m_out, 
    output logic sensor_r_out);



endmodule
