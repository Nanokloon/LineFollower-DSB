module robot
   (input logic clk,
    input logic reset,

    input logic sensor_l_in,
    input logic sensor_m_in,
    input logic sensor_r_in,

    output logic motor_l_pwm,
    output logic motor_r_pwm);



endmodule
